`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:13:56 04/30/2016 
// Design Name: 
// Module Name:    Video_Port 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Video_Port(
    input [7:0] DATA_IN,
    input STROBE,
    input HREF,
    input PCLK,
    input VSYNC,
    output XCLK,
    output RESET,
    output PWDN,
    output [7:0] DATA_OUT
    );


endmodule
