`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:13:50 04/30/2016 
// Design Name: 
// Module Name:    SCCB_Master_Unit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SCCB_Master_Unit(
    output IF_CLK,
    inout IF_DATA,
    input [6:0] ADDR,
    input [7:0] DATA_IN,
    output [7:0] DATA_OUT,
    input SEL,
    input RW
    );


endmodule
